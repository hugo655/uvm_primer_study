package my_pkg;
 import uvm_pkg::*;
 `include "uvm_macros.svh"


`include "dice_roller.svh"
`include "averager.svh"
`include "histogram.svh"
`include "main_test.svh"

endpackage
