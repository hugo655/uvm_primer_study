package my_pkg;
 import uvm_pkg::*;
 `include "uvm_macros.svh"


`include "main_test.svh"

endpackage
