class lion extends animal;


  function new(int a, string s);
    super.new(.a(a),.name(s));
  endfunction
  
  function void make_sound();
    $display("Lion makes ROAAAH");
  endfunction
endclass
