`include "verilog_dut/one_cycle_add_and_xor.sv"
`include "verilog_dut/three_cycle_mult.sv"
`include "verilog_dut/tiny_alu.sv"
