class lion_cage;
  static lion cage[$]; // Queue: an "array" which you don't know the length yet
endclass
