module top;

import uvm_pkg::*;
`include "uvm_macros.svh"

import my_pkg::*;

initial begin
  run_test();
end
endmodule : top
